// ed_sim_mem.v

// Generated using ACDS version 22.2 81

`timescale 1 ps / 1 ps
module ed_sim_mem (
		input  wire [0:0]  mem_ck,      // mem.mem_ck,      CK clock
		input  wire [0:0]  mem_ck_n,    //    .mem_ck_n,    CK clock (negative leg)
		input  wire [16:0] mem_a,       //    .mem_a,       Address
		input  wire [0:0]  mem_act_n,   //    .mem_act_n,   Activation command
		input  wire [1:0]  mem_ba,      //    .mem_ba,      Bank address
		input  wire [1:0]  mem_bg,      //    .mem_bg,      Bank group
		input  wire [0:0]  mem_cke,     //    .mem_cke,     Clock enable
		input  wire [0:0]  mem_cs_n,    //    .mem_cs_n,    Chip select
		input  wire [0:0]  mem_odt,     //    .mem_odt,     On-die termination
		input  wire [0:0]  mem_reset_n, //    .mem_reset_n, Asynchronous reset
		input  wire [0:0]  mem_par,     //    .mem_par,     Command and address parity
		output wire [0:0]  mem_alert_n, //    .mem_alert_n, Alert flag
		inout  wire [8:0]  mem_dqs,     //    .mem_dqs,     Data strobe
		inout  wire [8:0]  mem_dqs_n,   //    .mem_dqs_n,   Data strobe (negative leg)
		inout  wire [71:0] mem_dq,      //    .mem_dq,      Read/write data
		inout  wire [8:0]  mem_dbi_n    //    .mem_dbi_n,   Acts as either the data bus inversion pin, or the data mask pin, depending on configuration.
	);

	ed_sim_mem_altera_emif_mem_model_191_jkh6tsy mem (
		.mem_ck      (mem_ck),      //   input,   width = 1, mem.mem_ck
		.mem_ck_n    (mem_ck_n),    //   input,   width = 1,    .mem_ck_n
		.mem_a       (mem_a),       //   input,  width = 17,    .mem_a
		.mem_act_n   (mem_act_n),   //   input,   width = 1,    .mem_act_n
		.mem_ba      (mem_ba),      //   input,   width = 2,    .mem_ba
		.mem_bg      (mem_bg),      //   input,   width = 2,    .mem_bg
		.mem_cke     (mem_cke),     //   input,   width = 1,    .mem_cke
		.mem_cs_n    (mem_cs_n),    //   input,   width = 1,    .mem_cs_n
		.mem_odt     (mem_odt),     //   input,   width = 1,    .mem_odt
		.mem_reset_n (mem_reset_n), //   input,   width = 1,    .mem_reset_n
		.mem_par     (mem_par),     //   input,   width = 1,    .mem_par
		.mem_alert_n (mem_alert_n), //  output,   width = 1,    .mem_alert_n
		.mem_dqs     (mem_dqs),     //   inout,   width = 9,    .mem_dqs
		.mem_dqs_n   (mem_dqs_n),   //   inout,   width = 9,    .mem_dqs_n
		.mem_dq      (mem_dq),      //   inout,  width = 72,    .mem_dq
		.mem_dbi_n   (mem_dbi_n)    //   inout,   width = 9,    .mem_dbi_n
	);

endmodule
